library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity promDecimals is
    Port ( 
            addr      : in std_logic_vector(3 downto 0);
            keyCode   : in std_logic_vector(7 downto 0);
            M         : out std_logic_vector(31 downto 0)
    );
end promDecimals;

architecture Behavioral of promDecimals is

type memory_type is array (0 to 15) of std_logic_vector(31 downto 0);
    
---------------------------------------------------------------------------------
signal data_0 : memory_type :=(
							"11111111111111111111111111111111",
							"00000000000000000000000000000000",
							"00000000000000000000000111100000",
							"00000000000000000000011101110000",
							"00000000000000000000111000011100",
							"00000000000000000000111000011100",
							"00000000000000000000111000011100",
							"00000000000000000000111000011100",
							"00000000000000000000111000011100",
							"00000000000000000000111000011100",
							"00000000000000000000111000011100",
							"00000000000000000000011100011100",
							"00000000000000000000001110111000",
							"00000000000000000000000111000000",
							"00000000000000000000000000000000",
							"00000000000000000000000000000000"
							);
---------------------------------------------------------------------------------
signal data_1 : memory_type :=(
							"11111111111111111111111111111111",
							"00000000000000000000000000000000",
							"00000000000000000000000011111000",
							"00000000000000000000000110111000",
							"00000000000000000000011000111000",
							"00000000000000000000000000111000",
							"00000000000000000000000000111000",
							"00000000000000000000000000111000",
							"00000000000000000000000000111000",
							"00000000000000000000000000111000",
							"00000000000000000000000000111000",
							"00000000000000000000001111111111",
							"00000000000000000000000000000000",
							"00000000000000000000000000000000",
							"00000000000000000000000000000000",
							"00000000000000000000000000000000"
							);
---------------------------------------------------------------------------------
signal data_2 : memory_type :=(
							"11111111111111111111111111111111",
							"00000000000000000000000000000000",
							"00000000000000000000011111110000",
							"00000000000000000000111000111000",
							"00000000000000000001110000011100",
							"00000000000000000000000000011100",
							"00000000000000000000000000011100",
							"00000000000000000000000001110000",
							"00000000000000000000000011100000",
							"00000000000000000000000111000000",
							"00000000000000000000001110000000",
							"00000000000000000000001110000000",
							"00000000000000000000011111111100",
							"00000000000000000000111111111100",
							"00000000000000000000000000000000",
							"00000000000000000000000000000000"
							);
---------------------------------------------------------------------------------
signal data_3 : memory_type :=(
							"11111111111111111111111111111111",
							"00000000000000000000000000000000",
							"00000000000000000000111111110000",
							"00000000000000000001110000011100",
							"00000000000000000011100000011100",
							"00000000000000000000000000011100",
							"00000000000000000000000000111000",
							"00000000000000000000111111110000",
							"00000000000000000000000000111000",
							"00000000000000000000000000011100",
							"00000000000000000011100000011100",
							"00000000000000000001110000111000",
							"00000000000000000000011111110000",
							"00000000000000000000000000000000",
							"00000000000000000000000000000000",
							"00000000000000000000000000000000"
							);
---------------------------------------------------------------------------------
signal data_4 : memory_type :=(
							"11111111111111111111111111111111",
							"00000000000000000000000000000000",
							"00000000000000000000000011111000",
							"00000000000000000000000110111000",
							"00000000000000000000011000111000",
							"00000000000000000000110000111000",
							"00000000000000000001100000111000",
							"00000000000000000011000000111000",
							"00000000000000000111111111111000",
							"00000000000000000000000000111000",
							"00000000000000000000000000111000",
							"00000000000000000000000000111000",
							"00000000000000000000000000111000",
							"00000000000000000000001111111111",
							"00000000000000000000000000000000",
							"00000000000000000000000000000000"
							);
---------------------------------------------------------------------------------
signal data_5 : memory_type :=(
							"11111111111111111111111111111111",
							"00000000000000001111111111111000",
							"00000000000000001111111111111000",
							"00000000000000001110000000000000",
							"00000000000000001110000000000000",
							"00000000000000001110000000000000",
							"00000000000000001110000000000000",
							"00000000000000000111111000000000",
							"00000000000000000000001111000000",
							"00000000000000000000000001110000",
							"00000000000000000000000000111000",
							"00000000000000011100000001110000",
							"00000000000000011100000011100000",
							"00000000000000000111111110000000",
							"00000000000000000001111100000000",
							"00000000000000000000000000000000"
							);
---------------------------------------------------------------------------------
signal data_6 : memory_type :=(
							"11111111111111111111111111111111",
							"00000000000000000000000000000000",
							"00000000000000000000111111110000",
							"00000000000000000001110000000000",
							"00000000000000000011100000000000",
							"00000000000000000011100000000000",
							"00000000000000000011100000000000",
							"00000000000000000011111111110000",
							"00000000000000000011100000111000",
							"00000000000000000011100000011100",
							"00000000000000000011100000011100",
							"00000000000000000001110000111000",
							"00000000000000000000011111110000",
							"00000000000000000000000000000000",
							"00000000000000000000000000000000",
							"00000000000000000000000000000000"
							);
---------------------------------------------------------------------------------
signal data_7 : memory_type :=(
							"11111111111111111111111111111111",
							"00000000000000000000000000000000",
							"00000000000000000000000000000000",
							"00000000000000000011111111111100",
							"00000000000000000011111111111100",
							"00000000000000000000000000011100",
							"00000000000000000000000000011100",
							"00000000000000000000000001110000",
							"00000000000000000000000011100000",
							"00000000000000000000000111000000",
							"00000000000000000000001110000000",
							"00000000000000000000011100000000",
							"00000000000000000000111000000000",
							"00000000000000000000111000000000",
							"00000000000000000000000000000000",
							"00000000000000000000000000000000"
							);
---------------------------------------------------------------------------------
signal data_8 : memory_type :=(
							"11111111111111111111111111111111",
							"00000000000000000000000000000000",
							"00000000000000000000111111110000",
							"00000000000000000001110000011000",
							"00000000000000000011100000011100",
							"00000000000000000011100000011100",
							"00000000000000000011100000011100",
							"00000000000000000011111111110000",
							"00000000000000000011100000111000",
							"00000000000000000011100000011100",
							"00000000000000000011100000011100",
							"00000000000000000001110000111000",
							"00000000000000000000011111110000",
							"00000000000000000000000000000000",
							"00000000000000000000000000000000",
							"00000000000000000000000000000000"
							);
---------------------------------------------------------------------------------
signal data_9 : memory_type :=(
							"11111111111111111111111111111111",
							"00000000000000000000000000000000",
							"00000000000000000111111111111000",
							"00000000000000000111000000111000",
							"00000000000000000111000000111000",
							"00000000000000000111000000111000",
							"00000000000000000111000000111000",
							"00000000000000000111000000111000",
							"00000000000000000111111111111000",
							"00000000000000000000000000111000",
							"00000000000000000000000000111000",
							"00000000000000000000000000111000",
							"00000000000000000000000000111000",
							"00000000000000000000000000111000",
							"00000000000000000000000000111000",
							"00000000000000000000000000000000"
							);
---------------------------------------------------------------------------------
signal data_s : memory_type :=(
							"11111111111111111111111111111111",
							"00000000000000000000000000000000",
							"00000000000000000000000000000000",
							"00000000000000111110000000000000",
							"00000000000000111110000000000000",
							"00000000000000111110000000000000",
							"00000000000000000000000000000000",
							"00000000000000000000000000000000",
							"00000000000000000000000000000000",
							"00000000000000111110000000000000",
							"00000000000000111110000000000000",
							"00000000000000111110000000000000",
							"00000000000000000000000000000000",
							"00000000000000000000000000000000",
							"00000000000000000000000000000000",
							"00000000000000000000000000000000"
							);
---------------------------------------------------------------------------------
signal data_black : memory_type :=(
							"11111111111111111111111111111111",
							"00000000000000000000000000000000",
							"00000000000000000000000000000000",
							"00000000000000000000000000000000",
							"00000000000000000000000000000000",
							"00000000000000000000000000000000",
							"00000000000000000000000000000000",
							"00000000000000000000000000000000",
							"00000000000000000000000000000000",
							"00000000000000000000000000000000",
							"00000000000000000000000000000000",
							"00000000000000000000000000000000",
							"00000000000000000000000000000000",
							"00000000000000000000000000000000",
							"00000000000000000000000000000000",
							"00000000000000000000000000000000"
							);
---------------------------------------------------------------------------------

begin

    process(keyCode, addr)
    begin
        case keyCode is
           when "00000000" =>
              M <= data_0(to_integer(unsigned(addr)));
           when "00000001" =>
              M <= data_1(to_integer(unsigned(addr)));
           when "00000010" =>
              M <= data_2(to_integer(unsigned(addr)));
           when "00000011" =>
              M <= data_3(to_integer(unsigned(addr)));
           when "00000100" =>
              M <= data_4(to_integer(unsigned(addr)));
           when "00000101" =>
              M <= data_5(to_integer(unsigned(addr)));
           when "00000110" =>
              M <= data_6(to_integer(unsigned(addr)));
           when "00000111" =>
              M <= data_7(to_integer(unsigned(addr)));
           when "00001000" =>
              M <= data_8(to_integer(unsigned(addr)));
           when "00001001" =>
              M <= data_9(to_integer(unsigned(addr)));
           when "00001010" =>
              M <= data_s(to_integer(unsigned(addr)));
           when others =>
              M <= data_black(to_integer(unsigned(addr)));
        end case;
    end process;

end Behavioral;
